module adder(
    input [31:0] a
    );
endmodule

module adder(
    input logic [31:0] a
    );
endmodule