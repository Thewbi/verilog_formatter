module imem(
    input wire [31:0] a,
    output wire [31:0] rd);

    wire [31:0] RAM[63:0];

    initial
        $readmemh("riscvtest.txt", RAM);

    assign rd = RAM[a[31:2]]; // word aligned
endmodule