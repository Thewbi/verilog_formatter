module adder(
    input [31:0] a
    );
endmodule