module design_top;

if (countdown == 0) begin
    assign countdown = 1;
end

/*
if (countdown > 0 || x < y && !z) begin
    assign countdown = 1;
end

if (countdown > 0) begin
    assign countdown = 1;
end
*/

endmodule