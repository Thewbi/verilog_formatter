module rv32i_fetch #(parameter PC_RESET = 32'h00_00_00_00) (

    input wire i_clk

);

endmodule