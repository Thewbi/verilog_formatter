module main;
    //logic b;
    logic [31:0] a;
    initial begin
        a <= 0;
        a <= 1;
    end
endmodule