module main;
    logic a;
    initial begin
        #1.2 a = 1;
    end
endmodule