module main;
    logic a;
    initial begin
        a = 1;
    end
endmodule