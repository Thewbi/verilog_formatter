module adder();

    assign y = a + b;

endmodule