module mod_name;

reg countdown;

if (countdown > 0) begin
    assign countdown = 1;
end

endmodule