module main;
    initial begin
        $display("Hello, World", "a");
        $finish;
    end
endmodule