module top;

    initial begin
        $display("test");
    end

endmodule