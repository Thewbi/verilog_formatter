// implicit data type
module adder(
    input [31:0] a
    );
endmodule

// // explicit data type
// module adder(
//     input integer [31:0] a
//     );
// endmodule