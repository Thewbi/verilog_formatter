module testbench();
    adder dut(a, b, y);
endmodule
