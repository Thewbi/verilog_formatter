module wishbone_master (
//    input           i_reset,
//    input           i_cmd_stb,
    input   [33:0]	i_cmd_word
//    output  reg	    o_cmd_busy,
//    output          o_rsp_stb,
//    output          o_rsp_word
);

endmodule