module testbench();
    logic [31:0] a;
endmodule