module main;
    logic a;
    initial begin
        a <= 0;
        a <= 1;
    end
endmodule