module design_top;
    if (countdown > 0) begin
        assign countdown = 1;
    end
endmodule